LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY work;

ENTITY display IS
	PORT
	(
    	S0 :  IN  STD_LOGIC;
    	S1 :  IN  STD_LOGIC;
    	S2 :  IN  STD_LOGIC;
    	S3 :  IN  STD_LOGIC;
    	p0 :  OUT  STD_LOGIC;
    	p1 :  OUT  STD_LOGIC;
    	p2 :  OUT  STD_LOGIC;
    	p3 :  OUT  STD_LOGIC;
    	p4 :  OUT  STD_LOGIC;
    	p5 :  OUT  STD_LOGIC;
    	p6 :  OUT  STD_LOGIC
	);
END display;

ARCHITECTURE bdf_type OF display IS

SIGNAL	SYNTHESIZED_WIRE_123 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_124 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_125 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_126 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_127 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_128 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_129 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_130 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_131 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_132 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_133 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_134 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_135 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_136 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_137 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_138 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_139 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_140 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_141 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_142 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_119 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_120 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_121 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_122 :  STD_LOGIC;


BEGIN



SYNTHESIZED_WIRE_129 <= SYNTHESIZED_WIRE_123 AND SYNTHESIZED_WIRE_124 AND SYNTHESIZED_WIRE_125 AND SYNTHESIZED_WIRE_126;


SYNTHESIZED_WIRE_139 <= S0 AND SYNTHESIZED_WIRE_124 AND SYNTHESIZED_WIRE_125 AND SYNTHESIZED_WIRE_126;


SYNTHESIZED_WIRE_135 <= SYNTHESIZED_WIRE_123 AND S1 AND SYNTHESIZED_WIRE_125 AND S3;


SYNTHESIZED_WIRE_142 <= S0 AND S1 AND SYNTHESIZED_WIRE_125 AND S3;


SYNTHESIZED_WIRE_137 <= SYNTHESIZED_WIRE_123 AND SYNTHESIZED_WIRE_124 AND S2 AND S3;


SYNTHESIZED_WIRE_141 <= S0 AND SYNTHESIZED_WIRE_124 AND S2 AND S3;


SYNTHESIZED_WIRE_136 <= SYNTHESIZED_WIRE_123 AND S1 AND S2 AND S3;


SYNTHESIZED_WIRE_138 <= S0 AND S1 AND S2 AND S3;


SYNTHESIZED_WIRE_128 <= SYNTHESIZED_WIRE_123 AND S1 AND SYNTHESIZED_WIRE_125 AND SYNTHESIZED_WIRE_126;


SYNTHESIZED_WIRE_127 <= S0 AND S1 AND SYNTHESIZED_WIRE_125 AND SYNTHESIZED_WIRE_126;


SYNTHESIZED_WIRE_140 <= SYNTHESIZED_WIRE_123 AND SYNTHESIZED_WIRE_124 AND S2 AND SYNTHESIZED_WIRE_126;


SYNTHESIZED_WIRE_132 <= S0 AND SYNTHESIZED_WIRE_124 AND S2 AND SYNTHESIZED_WIRE_126;


SYNTHESIZED_WIRE_131 <= SYNTHESIZED_WIRE_123 AND S1 AND S2 AND SYNTHESIZED_WIRE_126;


SYNTHESIZED_WIRE_130 <= S0 AND S1 AND S2 AND SYNTHESIZED_WIRE_126;


SYNTHESIZED_WIRE_134 <= SYNTHESIZED_WIRE_123 AND SYNTHESIZED_WIRE_124 AND SYNTHESIZED_WIRE_125 AND S3;


SYNTHESIZED_WIRE_133 <= S0 AND SYNTHESIZED_WIRE_124 AND SYNTHESIZED_WIRE_125 AND S3;


p0 <= NOT(SYNTHESIZED_WIRE_32);



p1 <= NOT(SYNTHESIZED_WIRE_33);



p6 <= NOT(SYNTHESIZED_WIRE_34);



SYNTHESIZED_WIRE_123 <= NOT(S0);



SYNTHESIZED_WIRE_32 <= SYNTHESIZED_WIRE_127 OR SYNTHESIZED_WIRE_128 OR SYNTHESIZED_WIRE_129 OR SYNTHESIZED_WIRE_130 OR SYNTHESIZED_WIRE_131 OR SYNTHESIZED_WIRE_132 OR SYNTHESIZED_WIRE_133 OR SYNTHESIZED_WIRE_134 OR SYNTHESIZED_WIRE_135 OR SYNTHESIZED_WIRE_136 OR SYNTHESIZED_WIRE_137 OR SYNTHESIZED_WIRE_138;


SYNTHESIZED_WIRE_33 <= SYNTHESIZED_WIRE_128 OR SYNTHESIZED_WIRE_139 OR SYNTHESIZED_WIRE_129 OR SYNTHESIZED_WIRE_130 OR SYNTHESIZED_WIRE_140 OR SYNTHESIZED_WIRE_127 OR SYNTHESIZED_WIRE_133 OR SYNTHESIZED_WIRE_134 OR SYNTHESIZED_WIRE_135 OR SYNTHESIZED_WIRE_141 OR SYNTHESIZED_WIRE_141 OR SYNTHESIZED_WIRE_141;


SYNTHESIZED_WIRE_119 <= SYNTHESIZED_WIRE_127 OR SYNTHESIZED_WIRE_139 OR SYNTHESIZED_WIRE_129 OR SYNTHESIZED_WIRE_131 OR SYNTHESIZED_WIRE_132 OR SYNTHESIZED_WIRE_140 OR SYNTHESIZED_WIRE_134 OR SYNTHESIZED_WIRE_130 OR SYNTHESIZED_WIRE_133 OR SYNTHESIZED_WIRE_142 OR SYNTHESIZED_WIRE_135 OR SYNTHESIZED_WIRE_141;


SYNTHESIZED_WIRE_120 <= SYNTHESIZED_WIRE_127 OR SYNTHESIZED_WIRE_128 OR SYNTHESIZED_WIRE_129 OR SYNTHESIZED_WIRE_134 OR SYNTHESIZED_WIRE_131 OR SYNTHESIZED_WIRE_132 OR SYNTHESIZED_WIRE_142 OR SYNTHESIZED_WIRE_133 OR SYNTHESIZED_WIRE_137 OR SYNTHESIZED_WIRE_136 OR SYNTHESIZED_WIRE_141 OR SYNTHESIZED_WIRE_136;


SYNTHESIZED_WIRE_121 <= SYNTHESIZED_WIRE_131 OR SYNTHESIZED_WIRE_128 OR SYNTHESIZED_WIRE_129 OR SYNTHESIZED_WIRE_142 OR SYNTHESIZED_WIRE_135 OR SYNTHESIZED_WIRE_134 OR SYNTHESIZED_WIRE_141 OR SYNTHESIZED_WIRE_137 OR SYNTHESIZED_WIRE_136 OR SYNTHESIZED_WIRE_138 OR SYNTHESIZED_WIRE_138 OR SYNTHESIZED_WIRE_138;


SYNTHESIZED_WIRE_122 <= SYNTHESIZED_WIRE_132 OR SYNTHESIZED_WIRE_140 OR SYNTHESIZED_WIRE_129 OR SYNTHESIZED_WIRE_133 OR SYNTHESIZED_WIRE_134 OR SYNTHESIZED_WIRE_131 OR SYNTHESIZED_WIRE_142 OR SYNTHESIZED_WIRE_135 OR SYNTHESIZED_WIRE_137 OR SYNTHESIZED_WIRE_138 OR SYNTHESIZED_WIRE_136 OR SYNTHESIZED_WIRE_138;


SYNTHESIZED_WIRE_34 <= SYNTHESIZED_WIRE_140 OR SYNTHESIZED_WIRE_127 OR SYNTHESIZED_WIRE_128 OR SYNTHESIZED_WIRE_134 OR SYNTHESIZED_WIRE_131 OR SYNTHESIZED_WIRE_132 OR SYNTHESIZED_WIRE_135 OR SYNTHESIZED_WIRE_133 OR SYNTHESIZED_WIRE_142 OR SYNTHESIZED_WIRE_136 OR SYNTHESIZED_WIRE_141 OR SYNTHESIZED_WIRE_138;


SYNTHESIZED_WIRE_124 <= NOT(S1);



SYNTHESIZED_WIRE_125 <= NOT(S2);



SYNTHESIZED_WIRE_126 <= NOT(S3);



p2 <= NOT(SYNTHESIZED_WIRE_119);



p3 <= NOT(SYNTHESIZED_WIRE_120);



p4 <= NOT(SYNTHESIZED_WIRE_121);



p5 <= NOT(SYNTHESIZED_WIRE_122);



END bdf_type;